`timescale 1ns/1ps

module tb_cpu;
    // Signal declarations
    reg clk;                  // Clock signal
    reg reset;                // Reset signal
    wire [3:0] acc;           // Accumulator output from CPU module

    // Instantiate the CPU module under test (UUT)
    cpu uut (
        .clk(clk),
        .reset(reset),
        .acc(acc)
    );

    // Clock generation: 10 ns period (50 MHz)
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Test sequence
    initial begin
        // Enable GTKWave dump file generation
        $dumpfile("cpu_test.vcd");   // Specify the .vcd file name
        $dumpvars(0, tb_cpu);        // Record all variables in the tb_cpu module

        // Enhanced Monitor Statement for Readability
        $monitor("Time = %0dns | PC = %h | ACC (Accumulator) = %h | IR (Instruction) = %h | Operand = %b | Opcode = %b | R0 = %b | R1 = %b | ALU Output = %b",
                 $time, uut.PC, acc, uut.IR, uut.operand, uut.opcode, uut.R0, uut.R1, uut.alu_out);

        // Initialize the reset signal
        reset = 1;                     // Activate reset
        #10;
        reset = 0;                     // Release reset

        // Load instructions into memory from the "program.bin" file generated by the assembler
        $readmemb("program.bin", uut.memory);

        // Run the simulation for a sufficient time to observe instruction execution
        #400;

        // End simulation
        $finish;
    end
endmodule